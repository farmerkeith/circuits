* /home/guy/aProjects/circuits/regulator/regulatorTL431/regulatorTL431.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Sat 26 May 2018 19:11:32 AEST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
V1  Vin GND +13V 		
XQ1  Vg Vout Vin IRF4905		;Node Sequence Spec.<2,1,3>
R3  Vout GND 12		
R4  Vdiv GND 25K		
R2  Vout Vd 100K		
XD1  Vd GND Vdiv TL431		
R1  Vin Vg 500K		
R6  Vdiv Vout 103.37K		
Q1  Vg Vd Vdiv 2N3904		;Node Sequence Spec.<3,2,1>

*.include ../../ComponentModels/1n4148.spi
.include ../../ComponentModels/2n3904.spi
*.include ../../ComponentModels/ad822a.cir
.include ../../ComponentModels/irf4905.spi
.include ../../ComponentModels/tl431.spi
*.include ../../ComponentModels/1n4733.spi

.DC V1 0 20 0.1  
// DC analysis for 0 to 20 V in steps of 0.1V 

*.TRAN 1us 10ms
 // transient analysis for 10 ms in steps of 1 us (10,000 steps)
.control
run
plot vd vdiv vg title 'control voltages'
plot Vin Vout title 'input and output voltages'
plot Vin-Vout title 'drop out voltage'
plot Vin-Vout ylimit 0 0.05 title 'drop out voltage, expanded scale'
plot Vout ylimit 11.8 12.2 title 'output voltage, expanded scale'

.end
