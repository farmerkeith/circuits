* /home/guy/aProjects/circuits/currentShuntAmpDiscretesRes02/currentShuntAmpDiscretesRes02.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Wed 09 May 2018 11:25:14 AEST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
R4  Vout GND 10K		
Q1  Vc1 Vb1 VK 2N3906		
R5  Vc1 Vref 36K		
V1  VK GND +30V 		
I1  GND VA 1Amp		;Node Sequence Spec.<2,1>
R1  VK VA 4m		
R2  VA Ve1 63.65		
D1  Vref VK D1N4733		;Node Sequence Spec.<2,1>
R3  Vref GND 15K		
Q3  VC3 VB3 VE3 2N3906		
R6  VI3 VD2 8495.75		
R7  VD2 GND 15K		
D2  VD2 VK D1N4733		;Node Sequence Spec.<2,1>
R8  VK VE3 1		
R9  VB3 VI3 1		
R10  VC3 VI3 1		
R11  Vc1 Vb2 10m		
R12  Vb1 Vc1 10m		
Q2  Vout Vb2 Ve1 2N3906		

*.include ../ComponentModels/1n4148.spi
.include ../ComponentModels/2n3906.spi
*.include ../ComponentModels/irf4905.spi
.model D1N4733 D(Is=1.214f Rs=1.078 Ikf=0 N=1 Xti=3 Eg=1.11
+ Cjo=185p M=.3509 Vj=.75 Fc=.5  Bv=5.1 Ibv=.70507
+ Nbv=.74348 )
* Motorola pid=1N4733 case=DO-41

.DC I1 -0 8 0.01 // V1 20 40 10 
// DC analysis for 20, 30 and 40 Volts
//.DC I1 -0.5 8.5 0.1
// DC analysis from -0.5 to 8.5 Amps in steps of 0.1 Amp

*.TRAN 0.05us 10ms
 // transient analysis for 10 ms in steps of 0.1 us (10,000 steps)
.control
run
*plot Va Ve1 Vk
*plot (VA-VK)*25+2.693 Vout
*plot (VA-VK)*25+2.693-Vout
*plot VA VK  Vbase
*plot VK-Vref
*plot Ve1-Vc1 VA-Ve1 VA-Vc1 VK-Vc1
plot vout

.end
