* /home/guy/aProjects/circuits/currentShuntAmpDiscretes/currentShuntAmpDiscretes.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Sun 29 Apr 2018 15:15:38 AEST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
Q1  VC Vbase VA 2N3906		
R3  VC Vout 52.5K		
Q2  Vbase Vbase VK 2N3906		
R4  Vbase GND 280K		
R2  Net-_R2-Pad1_ VK 0		
V1  Net-_R2-Pad1_ GND +12V 		
R5  Vout GND 37.5K		
I1  GND VA 1Amp		;Node Sequence Spec.<2,1>
R1  VK VA 10m		

*.include ../ComponentModels/1n4148.spi
.include ../ComponentModels/2n3906.spi
*.include ../ComponentModels/irf4905.spi

.DC I1 -5 5 0.1
// DC analysis from 0 to 1 Amps in steps of 1 Amp
*.TRAN 0.05us 10ms
 // transient analysis for 10 ms in steps of 0.1 us (10,000 steps)
.control
run
plot VA VK  VC Vbase
plot (VA-VK)
plot (VA-VK)*50+2.5 Vout

.end
