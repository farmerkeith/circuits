* /home/guy/aProjects/circuits/MOSFETdiodeDiscretesHiV/MOSFETdiodeDiscretesHiV.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Sun 13 May 2018 09:48:43 AEST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
D1  VA Net-_D1-Pad1_ 1N4148		;Node Sequence Spec.<2,1>
D2  VK Net-_D2-Pad1_ 1N4148		;Node Sequence Spec.<2,1>
Q2  Vbase Vbase Net-_D1-Pad1_ 2N3906		
R2  Vbase VD 470K		
Q3  VG Vbase Net-_D2-Pad1_ 2N3906		
R3  VG VD 470K		
V1  VA GND 25V		
R1  Net-_R1-Pad1_ VK 10		
V2  Net-_R1-Pad1_ GND +40V 		
R4  VD GND 100K		
XQ1  VA VG VK IRF4905		
D3  VD VK 1N4742 		;Node Sequence Spec.<2,1>

.include ../ComponentModels/1n4148.spi
.include ../ComponentModels/2n3906.spi
.include ../ComponentModels/irf4905.spi
.include ../ComponentModels/1n4742.spi

.DC V1 25 45 1
*.TRAN 0.05us 10ms
 // transient analysis for 10 ms in steps of 0.1 us (10,000 steps)
*pulse (9.50V 11.5V 2ms 0 0 5ms 10ms 0) V1 for transient analysis
.control
run
plot VA VK  VG Vbase
plot VA-VK
plot VA-Vbase VK-Vbase VK-VG
plot -i(V1) i(V2)
plot VD VK-VD

.end
