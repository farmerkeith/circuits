* /home/guy/aProjects/circuits/regulator/regulatorOpAmp/regulatorOpAmp.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Sat 26 May 2018 13:35:21 AEST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
V1  Vin GND +13V 		
XU1  Vdiv Vref Vin GND Vg AD822A		;Node Sequence Spec.<3,2,8,4,1>
R2  Vout Vref 115K		
XQ1  Vg Vout Vin IRF4905		;Node Sequence Spec.<2,1,3>
R3  Vout GND 6		
D1  Vref GND 1N4148		;Node Sequence Spec.<2,1>
R4  Vdiv GND 5K		
R1  Vout Vdiv 115.28K		

.include ../../ComponentModels/1n4148.spi
*.include ../../ComponentModels/2n3906.spi
.include ../../ComponentModels/ad822a.cir
.include ../../ComponentModels/irf4905.spi
*.include ../../ComponentModels/1n4733.spi

.DC V1 0 20 0.1  
// DC analysis for 0 to 20 V in steps of 0.1V 

*.TRAN 1us 10ms
 // transient analysis for 10 ms in steps of 1 us (10,000 steps)
.control
run
plot Vin-Vg Vref*20 Vdiv*20 title 'control voltages'
plot Vin Vout title 'input and output voltages'
plot Vin-Vout title 'drop out voltage'
plot Vin-Vout ylimit 0 0.05 title 'drop out voltage, expanded scale'
plot Vout ylimit 11.8 12.2 title 'output voltage, expanded scale'

.end
