* /home/guy/aProjects/circuits/mainsControl/mains/mains.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Mon 21 May 2018 21:15:34 AEST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
V1  Net-_R2-Pad2_ GND sine 0 340V 50Hz		
L1  VP GND 50H		
L2  VS VS2 124mH 		
R1  Net-_R1-Pad1_ VR 1		
R2  VP Net-_R2-Pad2_ 0.01R		
D1  GND VS 2W01G		;Node Sequence Spec.<2,1>
D3  GND VS2 2W01G		;Node Sequence Spec.<2,1>
D2  VS Net-_D2-Pad1_ 2W01G		;Node Sequence Spec.<2,1>
D4  VS2 Net-_D2-Pad1_ 2W01G		;Node Sequence Spec.<2,1>
C1  VR GND 10000uF		
V2  Net-_R1-Pad1_ GND DC 12V 		
R3  VR Net-_D2-Pad1_ 0.5		

.include ../../ComponentModels/2w01g.spi
K L1 L2 1
.TRAN 0.0001 0.1
.control
run
plot VP VS
plot i(v1)
plot vs vs2 vr
plot i(v2)
.end

.end
