* model from http://users.skynet.be/hugocoolens/spice/transist/bc547b.htm
*DATABOOK PHILIPS
.MODEL BC547B  NPN (BF=530 NE=1.3 ISE=9.72F IKF=80M IS=20F VAF=50V
+      BR=10 NC=2 ISC=47P IKR=12M VAR=10
+      RB=280 RE=1 RC=40 TR=.3U
+      CJE=12P VJE=.48 MJE=0.5 CJC=6P VJC=.7 MJC=.33 TF=.5N)
