* /home/guy/aProjects/circuits/currentShuntAmpDiscretesRes01/currentShuntAmpDiscretesRes01.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Tue 01 May 2018 23:48:40 AEST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
Q1  VC Vbase Net-_Q1-Pad3_ 2N3906		
R4  VC Vout 52.5K		
Q2  Vbase Vbase Net-_Q2-Pad3_ 2N3906		
R5  Vbase GND 240K		
V1  VK GND +12V 		
R6  Vout GND 37.5K		
I1  GND VA 1Amp		;Node Sequence Spec.<2,1>
R1  VK VA 10m		
R2  VA Net-_Q1-Pad3_ 1K		
R3  VK Net-_Q2-Pad3_ 1K		

*.include ../ComponentModels/1n4148.spi
.include ../ComponentModels/2n3906.spi
*.include ../ComponentModels/irf4905.spi

.DC I1 -12 12 0.1
// DC analysis from 0 to 1 Amps in steps of 1 Amp
*.TRAN 0.05us 10ms
 // transient analysis for 10 ms in steps of 0.1 us (10,000 steps)
.control
run
plot VA VK  VC Vbase
plot (VA-VK)
plot (VA-VK)*23.5+2.15 Vout
plot (VA-VK)*23.5+2.15-Vout

.end
