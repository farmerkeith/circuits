* /home/guy/aProjects/circuits/PWMdriver/voltageSources/voltageSources.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Fri 01 Jun 2018 18:17:19 AEST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
V2  VA 0 +12V		
R2  VSine 0 10K		
R1  VA 0 10K		
V3  VC 0 +5V		
R3  VC Net-_R3-Pad2_ 10K		
V4  Net-_R3-Pad2_ GND 0V		
R4  VPulse 0 10K		
V1  VSine 0 Vsine0VOffset17.1Vpeak50Hz1mSDelay0Damping0Phase		
V5  VPulse 0 Vpulse0VInit4.95Vpulsed2nSDelay0.2mSRise.2mSFall10.85mSWidth20mSPeriod0Phase		

.TRAN 0.1m 40m
.control
run
plot VA VSine VC title 'DC and sine voltages'
plot VPulse title 'pulse voltage'
plot VA VSine VPulse VC title 'Waveforms'

.end
