*file bs250p.spi
*spice model for P-channel MOSFET BS250P with KH comments 11 May 2018
* obtained from http://ltwiki.org/index.php?title=Bs250
* model consists of 3 capacitors, 2 MOSFETs and 1 body diode

.SUBCKT BS250P 2 1 3 // G D S 
* 1=drain 2=gate 3=source
 Cgs 2 3 20.1E-12  // Cap 20.1 pF G S
 Cgd1 2 4 57.1E-12 // Cap 57.1 pF G 4
 Cgd2 1 4 5E-12    // Cap 5 pF    D 4
 M1 1 2 3 3 MOST1  // MOSFET D G S S 
 M2 4 2 1 3 MOST2  // MOSFET 4 G D S 
 D1 1 3 Dbody      // DIODE      D S (body diode)

.MODEL MOST1 PMOS(LEVEL=3 // MOSFET
 + VTO=-2.3 // zero bias threshold voltage
 + W=7.6m   // channel width? Not accepted by ngspice
 + L=2u     // channel length? Not accepted by ngspice
 + KP=10.33u 
 + RD=4.014 
 + RS=20m) 
.MODEL MOST2 PMOS( // MOSFET
 + VTO=2.43 // zero bias threshold voltage
 + W=7.6m   // channel width? Not accepted by ngspice
 + L=2u     // channel length? Not accepted by ngspice
 + KP=10.33u 
 + RS=20m) 
.MODEL Dbody D(    // Diode
 + CJO=53.22E-12 
 + VJ=0.5392 
 + M=0.3583 
 + IS=75.32E-15 
 + N=1.016 
 + RS=1.245 
 + TT=86.56n 
 + BV=45        // breakdown voltage
 + IBV=10u) 
.ENDS
