*Package Pin 1 : Cathode
*Package Pin 2 : Anode

*.SUBCKT MBR2045 2 1 
*
* The resistor R1 does not reflect 
* a physical device. Instead it
* improves modeling in the reverse 
* mode of operation.
*
*R1 1 2 5.827E+9 
*D1 1 2 1N4148
*
.MODEL MBR2045 D 
+ IS = 1.62944E-5
+ N = 1.906 
+ BV = 45 
+ IBV = 0.0001 
+ RS = 0.0003
+ CJO = 1E-9 // guess  
+ VJ = 0.869 
+ M = 0.03 
+ FC = 0.5 
+ TT = 3.48E-9 

*.ENDS
