Model from http://vlabs.iitb.ac.in/vlab/electrical/resources/bc547.txt
*BC547BP ZETEX Spice model     Last revision  4/90   General Purpose
*ZTX Si 500mW  45V 200mA 300MHz pkg:TO-92 1,2,3
.MODEL QBC547BP NPN(IS=1.8E-14 BF=400 NF=0.9955 VAF=80 IKF=0.14 ISE=5E-14 
+ NE=1.46 BR=35.5 NR=1.005 VAR=12.5 IKR=0.03 ISC=1.72E-13 NC=1.27 RB=0.56 
+ RE=0.6 RC=0.25 CJE=1.3E-11 TF=6.4E-10 CJC=4E-12 VJC=0.54 TR=5.072E-8 )
