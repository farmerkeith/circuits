* /home/guy/aProjects/circuits/diodeTest/diodeTest.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Mon 21 May 2018 14:45:42 AEST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
V1  Net-_D1-Pad2_ GND DC 0V		
D1  Net-_D1-Pad2_ Net-_D1-Pad1_ 2W01G		;Node Sequence Spec.<2,1>
V2  Net-_D1-Pad1_ GND DC 0V		

.include ../ComponentModels/2w01g.spi
.DC V1 0.63 1.6 0.01 
.control
run
plot i(v2)
plot log(i(v2))/log(10)
end

.end
