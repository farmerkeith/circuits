.model bc547 NPN BF=400 NE=1.3 ISE=10.3F IKF=50M IS=10F VAF=80 ikr=12m
       + BR=9.5 NC=2 VAR=10 RB=280 RE=1 RC=40 VJE=.48 tr=.3u tf=.5n
       +cje=12p vje=.48 mje=.5 cjc=6p vjc=.7 mjc=.33 isc=47p kf=2f
.model bc547b NPN BF=500 NE=1.3 ISE=9.72F IKF=80M IS=20F VAF=50 ikr=12m
       + BR=10 NC=2 VAR=10 RB=280 RE=1 RC=40 VJE=.48 tr=.3u tf=.5n
       +cje=12p vje=.48 mje=.5 cjc=6p vjc=.7 mjc=.33 isc=47p kf=2f
.model bc547c NPN BF=730 NE=1.4 ISE=29.5F IKF=80M IS=60F VAF=25 ikr=12m
       + BR=10 NC=2 VAR=10 RB=280 RE=1 RC=40 VJE=.48 tr=.3u tf=.5n
       +cje=12p vje=.48 mje=.5 cjc=6p vjc=.7 mjc=.33 isc=47.6p kf=2f
.model BC557 PNP BF=190 NE=1.5 ISE=12F IKF=90M IS=10F VAF=50 ikr=12m
       + nc=2 br=4 var=10 rb=280 re=1 rc=40 vje=.48 tf=.5n tr=.3u
       +cje=12p vje=.48 mje=.5 cjc=6p vjc=.7 mjc=.33 isc=47.6p kf=2f
.model BC557b PNP BF=335 NE=1.5 ISE=7.35F IKF=82M IS=10F VAF=40 ikr=12m
       + nc=2 br=4 var=10 rb=280 re=1 rc=40 vje=.48 tf=.5n tr=.3u
       +cje=12p vje=.48 mje=.5 cjc=6p vjc=.7 mjc=.33 isc=47.6p kf=2f
.model BC557c PNP BF=490 NE=1.5 ISE=12.4F IKF=78M IS=60F VAF=36 ikr=12m
       + nc=2 br=4 var=10 rb=280 re=1 rc=40 vje=.48 tf=.5n tr=.3u
       +cje=12p vje=.48 mje=.5 cjc=6p vjc=.7 mjc=.33 isc=47.6p kf=2f
