* /home/guy/aProjects/circuits/NGspice/Schmidt/Schmidt.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Mon 04 Jun 2018 21:55:56 AEST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
R1  Vout GND 10K		
V1  Net-_E1-Pad3_ GND +12V		
E1  Net-_E1-Pad1_ GND Net-_E1-Pad3_ GND VCVS0.5Gain		
V2  Net-_S1-Pad1_ GND +5V		
V3  Vin GND Vpulse0VInit12Vpulsed2nsDelay2msRise2msFall8msWidth20msPeriod0Phase		
S1  Net-_S1-Pad1_ Vout Vin Net-_E1-Pad1_ Schmidt0.5VHysteresis		

.TRAN 0.1m 40m
.control
run
plot Vin Vout title 'Waveforms'

.end
