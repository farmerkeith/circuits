* /home/guy/aProjects/circuits/currentShuntAmpOpAmpUniMOS/currentShuntAmpOpAmpUniMOS.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Sat 12 May 2018 08:52:43 AEST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
V1  VK GND +30V 		
I1  GND VA 1Amp		;Node Sequence Spec.<2,1>
R1  VK VA 4m		
XU1  Net-_R4-Pad2_ Ve VK Vneg Vb AD822A		;Node Sequence Spec.<3,2,8,4,1>
R2  VA Ve 100R		
R3  Vout GND 15.665K		
D1  Vneg VK D1N4733		;Node Sequence Spec.<2,1>
R6  Vneg GND 10K		
R4  VK Net-_R4-Pad2_ 16.8		
R5  Net-_R4-Pad2_ Vneg 50K		
XQ1  Vb Vout Ve BS250P		

*.include ../ComponentModels/1n4148.spi
.include ../ComponentModels/2n3906.spi
.include ../ComponentModels/ad822a.cir
.include ../ComponentModels/bs250p.spi
*.include ../ComponentModels/irf4905.spi
.model D1N4733 D(Is=1.214f Rs=1.078 Ikf=0 N=1 Xti=3 Eg=1.11
+ Cjo=185p M=.3509 Vj=.75 Fc=.5  Bv=5.1 Ibv=.70507
+ Nbv=.74348 )
* Motorola pid=1N4733 case=DO-41

*.MODEL BS250P VDMOS pchan Rg=160 VTO=-3.193 RS=2.041 RD=0.697
*.MODEL MBS250P PMOS(Rg=160 VTO=-3.193 RS=2.041 RD=0.697
*+ IS=2E-13 KP=0.277 Cjo=105p PB=1 LAMBDA=1.2E-2 RB=0.309
*+Rds=1.2E8 Cgdmax=57p Cgdmin=5p CGS=47p TT=86.56n BV=45 IBV=10u)

.DC I1 0 8 0.1  V1 20 40 10 
*.DC I1 -0.1 0.8 0.01  
// DC analysis for 20, 30 and 40 Volts
//.DC I1 -0.5 8.5 0.1
// DC analysis from -0.5 to 8.5 Amps in steps of 0.1 Amp

*.TRAN 0.05us 10ms
 // transient analysis for 10 ms in steps of 0.1 us (10,000 steps)
.control
run
*plot Va Ve1 Vk
*plot (VA-VK)*25+2.693 Vout
*plot (VA-VK)*25+2.693-Vout
*plot VA VK  Vbase
*plot VK-Vref
*plot Ve1-Vc1 VA-Ve1 VA-Vc1 VK-Vc1
plot vout
plot vout-i(v1)*5/8 // voltage error
plot vout*8/5-i(v1) // ccurrent error
*plot i1

.end
