* /home/guy/aProjects/circuits/MOSFETdiode/MOSFETdiodeDiscretesHiV/MOSFETdiodeDiscretesHiV.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Fri 25 May 2018 22:32:00 AEST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
D1  VA Net-_D1-Pad1_ 1N4148		;Node Sequence Spec.<2,1>
D2  VK Net-_D2-Pad1_ 1N4148		;Node Sequence Spec.<2,1>
Q2  Vbase Vbase Net-_D1-Pad1_ 2N3906		
R2  Vbase VD 47K		
Q3  VG Vbase Net-_D2-Pad1_ 2N3906		
R3  VG VD 47K		
V1  VA GND pulse (25V 40V 2ms 0 0 5ms 10ms 0) //  25V // 		
R1  Net-_R1-Pad1_ VK 10		
V2  Net-_R1-Pad1_ GND +30V 		
R4  VD GND 27K		
XQ1  VG VA VK IRF4905		;Node Sequence Spec.<2,1,3>
D3  VD VK 1N4742 		;Node Sequence Spec.<2,1>

.include ../../ComponentModels/1n4148.spi
.include ../../ComponentModels/2n3906.spi
.include ../../ComponentModels/irf4905.spi
.include ../../ComponentModels/1n4742.spi

*.DC V1 -1 45 1 // DC analysis
.TRAN 100us 10ms
 // transient analysis for 10 ms in steps of 100 us (10,000 steps)
.control
run
plot VA VK  VG Vbase title "applied voltages"
plot VA-VK title "Forward Voltage"
plot VA-Vbase VK-Vbase VK-VG title "control voltages"
plot -i(V1) i(V2) title "currents"
plot VD VK-VD title "Zener offset"

.end
