* /home/guy/aProjects/circuits/PWMdriver/switchChangeover/switchChangeover.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Mon 04 Jun 2018 17:02:51 AEST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
V2  IN GND pulse 0V 5V 2ns 3us 3us 7us 20us  		
V1  Net-_S1-Pad2_ GND 12V 		
C1  OUT GND 10nF		
R1  OUT Net-_R1-Pad2_ 15		
R2  OUT Net-_R2-Pad2_ 15		
S1  Net-_R1-Pad2_ Net-_S1-Pad2_ IN GND SwitchNO		
S2  GND Net-_R2-Pad2_ IN GND SwitchNC		

.tran 5us 41us
.control 
run
plot in out  title 'Switching action'

.end
