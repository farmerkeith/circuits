* /home/guy/aProjects/circuits/PWMdriver/voltageSources/voltageSources.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Thu 31 May 2018 23:26:08 AEST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
V2  VA 0 +12V		
R2  VB 0 10K		
R1  VA 0 10K		
V3  VC 0 +5V		
R3  VC Net-_R3-Pad2_ 10K		
V1  VB 0 Vsine0VOffset17.1Vpeak50Hz1mSDelay0Damping0Phase		
V4  Net-_R3-Pad2_ GND 0V		

.TRAN 0.1m 40m
.control
run
plot VA VB VC title 'voltages'

.end
